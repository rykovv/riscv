module alu #(
  parameter WORDSIZE = 64
) (
  input [WORDSIZE-1:0] A, B,
  input [3:0] CTL,
  output z,
  output [WORDSIZE-1:0] R
);



endmodule
