`include "riscv.v"

module riscv_tb();
  reg clk;

endmodule
